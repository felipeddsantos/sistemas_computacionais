//Sistemas Computacionais - Unidade Lógica Aritmética (Somador 16)
//Felipe Daniel Dias dos Santos - 11711ECP004
//Graduação em Engenharia de Computação - Faculdade de Engenharia Elétrica - Universidade Federal de Uberlândia

CHIP Add16{

    IN a[16], b[16];
    OUT out[16];

    PARTS:

        HalfAdder(a = a[0], b = b[0], sum = out[0], carry = out1);
        FullAdder(a = a[1], b = b[1], c = out1, sum = out[1], carry = out2);
        FullAdder(a = a[2], b = b[2], c = out2, sum = out[2], carry = out3);
        FullAdder(a = a[3], b = b[3], c = out3, sum = out[3], carry = out4);
        FullAdder(a = a[4], b = b[4], c = out4, sum = out[4], carry = out5);
        FullAdder(a = a[5], b = b[5], c = out5, sum = out[5], carry = out6);
        FullAdder(a = a[6], b = b[6], c = out6, sum = out[6], carry = out7);
        FullAdder(a = a[7], b = b[7], c = out7, sum = out[7], carry = out8);
        FullAdder(a = a[8], b = b[8], c = out8, sum = out[8], carry = out9);
        FullAdder(a = a[9], b = b[9], c = out9, sum = out[9], carry = out10);
        FullAdder(a = a[10], b = b[10], c = out10, sum = out[10], carry = out11);
        FullAdder(a = a[11], b = b[11], c = out11, sum = out[11], carry = out12);
        FullAdder(a = a[12], b = b[12], c = out12, sum = out[12], carry = out13);
        FullAdder(a = a[13], b = b[13], c = out13, sum = out[13], carry = out14);
        FullAdder(a = a[14], b = b[14], c = out14, sum = out[14], carry = out15);
        FullAdder(a = a[15], b = b[15], c = out15, sum = out[15], carry = out16);
}                       
